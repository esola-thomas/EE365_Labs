library ieee;
use ieee.std_logic_1164.all;

package values is
	constant N: integer :=4;	-- must not be more than 6 for the DE0_Nano board	
	constant upper: integer :=13;	-- must not be more than 6 for the DE0_Nano board	
	constant lower: integer :=2;	-- must not be more than 6 for the DE0_Nano board		
end package values;