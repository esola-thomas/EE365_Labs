-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version
-- Created on Wed Sep 28 22:01:38 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY StateMachine_Rotary_Encoder IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        A : IN STD_LOGIC := '0';
        B : IN STD_LOGIC := '0';
        Add : OUT STD_LOGIC;
        Subtract : OUT STD_LOGIC
    );
END StateMachine_Rotary_Encoder;

ARCHITECTURE BEHAVIOR OF StateMachine_Rotary_Encoder IS
    TYPE type_fstate IS (CarStartsExit,CarStartsEnter,CarHalfWayIn,Load,CarHalfWayOut,In75,CarIn,Out75,CarOut);
    SIGNAL fstate : type_fstate := Load;
    SIGNAL reg_fstate : type_fstate := Load;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,A,B)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Load;
            Add <= '0';
            Subtract <= '0';
        ELSE
            Add <= '0';
            Subtract <= '0';
            CASE fstate IS
                WHEN CarStartsExit =>
                    IF (((A = '1') AND (B = '1'))) THEN
                        reg_fstate <= Load;
                    ELSIF (((A = '0') AND (B = '0'))) THEN
                        reg_fstate <= CarHalfWayOut;
                    ELSE
                        reg_fstate <= CarStartsExit;
                    END IF;
                WHEN CarStartsEnter =>
                    IF (((A = '1') AND (B = '1'))) THEN
                        reg_fstate <= Load;
                    ELSIF (((A = '0') AND (B = '0'))) THEN
                        reg_fstate <= CarHalfWayIn;
                    ELSE
                        reg_fstate <= CarStartsEnter;
                    END IF;
                WHEN CarHalfWayIn =>
                    IF (((A = '0') AND (B = '1'))) THEN
                        reg_fstate <= CarStartsEnter;
                    ELSIF (((A = '1') AND (B = '0'))) THEN
                        reg_fstate <= In75;
                    ELSE
                        reg_fstate <= CarHalfWayIn;
                    END IF;
                WHEN Load =>
                    IF (((A = '0') AND (B = '1'))) THEN
                        reg_fstate <= CarStartsEnter;
                    ELSIF (((A = '1') AND (B = '0'))) THEN
                        reg_fstate <= CarStartsExit;
                    ELSE
                        reg_fstate <= Load;
                    END IF;

                    Add <= '0';

                    Subtract <= '0';
                WHEN CarHalfWayOut =>
                    IF (((A = '1') AND (B = '0'))) THEN
                        reg_fstate <= CarStartsExit;
                    ELSIF (((A = '0') AND (B = '1'))) THEN
                        reg_fstate <= Out75;
                    ELSE
                        reg_fstate <= CarHalfWayOut;
                    END IF;
                WHEN In75 =>
                    IF (((A = '1') AND (B = '1'))) THEN
                        reg_fstate <= CarIn;
                    ELSIF (((A = '0') AND (B = '0'))) THEN
                        reg_fstate <= CarHalfWayIn;
                    ELSE
                        reg_fstate <= In75;
                    END IF;
                WHEN CarIn =>
                    reg_fstate <= Load;

                    Add <= '1';
                WHEN Out75 =>
                    IF (((A = '0') AND (B = '0'))) THEN
                        reg_fstate <= CarHalfWayOut;
                    ELSIF (((A = '1') AND (B = '1'))) THEN
                        reg_fstate <= CarOut;
                    ELSE
                        reg_fstate <= Out75;
                    END IF;
                WHEN CarOut =>
                    reg_fstate <= Load;

                    Subtract <= '1';
                WHEN OTHERS => 
                    Add <= '0';
                    Subtract <= '0';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
