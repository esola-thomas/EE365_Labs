-- Copyright (C) 2022  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 21.1.1 Build 850 06/23/2022 SJ Lite Edition
-- Created on Sat Oct  1 13:45:47 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY StateMachine_Rotary_Encoder IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        A : IN STD_LOGIC := '0';
        B : IN STD_LOGIC := '0';
        max : IN STD_LOGIC := '0';
        min : IN STD_LOGIC := '0';
        en : OUT STD_LOGIC;
        up : OUT STD_LOGIC;
        clk_en : OUT STD_LOGIC
    );
END StateMachine_Rotary_Encoder;

ARCHITECTURE BEHAVIOR OF StateMachine_Rotary_Encoder IS
    TYPE type_fstate IS (CarStartsExit,CarStartsEnter,CarHalfWayIn,Load,CarHalfWayOut,In75,CarIn,Out75,CarOut);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,A,B,max,min)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Load;
            en <= '0';
            up <= '0';
            clk_en <= '0';
        ELSE
            en <= '0';
            up <= '0';
            clk_en <= '0';
            CASE fstate IS
                WHEN CarStartsExit =>
                    IF (((A = '1') AND (B = '1'))) THEN
                        reg_fstate <= Load;
                    ELSIF (((A = '0') AND (B = '0'))) THEN
                        reg_fstate <= CarHalfWayOut;
                    ELSE
                        reg_fstate <= CarStartsExit;
                    END IF;
                WHEN CarStartsEnter =>
                    IF (((A = '1') AND (B = '1'))) THEN
                        reg_fstate <= Load;
                    ELSIF (((A = '0') AND (B = '0'))) THEN
                        reg_fstate <= CarHalfWayIn;
                    ELSE
                        reg_fstate <= CarStartsEnter;
                    END IF;
                WHEN CarHalfWayIn =>
                    IF (((A = '0') AND (B = '1'))) THEN
                        reg_fstate <= CarStartsEnter;
                    ELSIF (((A = '1') AND (B = '0'))) THEN
                        reg_fstate <= In75;
                    ELSE
                        reg_fstate <= CarHalfWayIn;
                    END IF;
                WHEN Load =>
                    IF ((((A = '0') AND (B = '1')) AND (max = '0'))) THEN
                        reg_fstate <= CarStartsEnter;
                    ELSIF ((((A = '1') AND (B = '0')) AND (min = '0'))) THEN
                        reg_fstate <= CarStartsExit;
                    ELSE
                        reg_fstate <= Load;
                    END IF;

                    clk_en <= '0';

                    en <= '0';
                WHEN CarHalfWayOut =>
                    IF (((A = '1') AND (B = '0'))) THEN
                        reg_fstate <= CarStartsExit;
                    ELSIF (((A = '0') AND (B = '1'))) THEN
                        reg_fstate <= Out75;
                    ELSE
                        reg_fstate <= CarHalfWayOut;
                    END IF;
                WHEN In75 =>
                    IF (((A = '1') AND (B = '1'))) THEN
                        reg_fstate <= CarIn;
                    ELSIF (((A = '0') AND (B = '0'))) THEN
                        reg_fstate <= CarHalfWayIn;
                    ELSE
                        reg_fstate <= In75;
                    END IF;
                WHEN CarIn =>
                    reg_fstate <= Load;

                    clk_en <= '1';

                    up <= '1';

                    en <= '1';
                WHEN Out75 =>
                    IF (((A = '0') AND (B = '0'))) THEN
                        reg_fstate <= CarHalfWayOut;
                    ELSIF (((A = '1') AND (B = '1'))) THEN
                        reg_fstate <= CarOut;
                    ELSE
                        reg_fstate <= Out75;
                    END IF;
                WHEN CarOut =>
                    reg_fstate <= Load;

                    clk_en <= '1';

                    up <= '0';

                    en <= '1';
                WHEN OTHERS => 
                    en <= '0';
                    up <= '0';
                    clk_en <= '0';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
