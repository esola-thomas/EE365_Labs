LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY keys IS
PORT ( CLOCK_50 : IN STD_LOGIC;
KEY : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
LED : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)); -- GREEN LEDs
END keys;
ARCHITECTURE Behavior OF keys IS
BEGIN
PROCESS (CLOCK_50)
BEGIN
IF(RISING_EDGE(CLOCK_50)) THEN
LED <= KEY;
END IF;
END PROCESS;
END Behavior;
